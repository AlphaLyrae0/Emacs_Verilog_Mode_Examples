module sub2 (
    interface if_int, // Generic Interface
    interface if_o    // Generic Interface
);

endmodule