module top 
(
    /*AUTOINPUT*/

    /*AUTOOUTPUT*/

);

    /*AUTOWIRE*/

    /* sub1 AUTO_TEMPLATE (
        .sig_a (a_top[]),
        .sig_b (b_top[]),
        .sig_c (c_top[][]),
        .sig_d (d_top[][]),
        .sig_e (e_top[]),
        .sig_f (f_top[]),
        .sig_g (g_top[][]),
        .sig_h (h_top[][]),
    ) */
    sub1    s1
    ( /*AUTOINST*/);

    /* sub2 AUTO_TEMPLATE (
        .sig_e (e_top[]),
        .sig_f (f_top[]),
        .sig_g (g_top[][]),
        .sig_h (h_top[][]),
        .sig_i (i_top[]),
        .sig_j (j_top[]),
        .sig_k (k_top[][]),
        .sig_l (l_top[][]),
    ) */
    sub2    s2
    (
        /*AUTOINST*/);

endmodule
// Local Variables:
// verilog-library-flags:("-y ./sub")
// verilog-auto-inst-column:24  ;; Min. 24?
// indent-tabs-mode:nil
// End:


// verilog-auto-inst-dot-name:t
// verilog-auto-inst-vector:nil
