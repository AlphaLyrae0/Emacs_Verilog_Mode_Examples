module top import my_pkg::*;
(
    /*AUTOINPUT*/

    /*AUTOOUTPUT*/

);

    /*AUTOWIRE*/

    sub1    s1
    ( /*AUTOINST*/);

    sub2    s2
    ( /*AUTOINST*/);

endmodule
// Local Variables:
// verilog-library-flags:("-y ./sub")
// verilog-auto-inst-column:24
// verilog-typedef-regexp:"_t$"
// indent-tabs-mode:nil
// End:

// verilog-typedef-regexp:"\\(_t$\\|_st$\\|_e$\\|^t_\\)"
// verilog-auto-inst-dot-name:t
// verilog-auto-inst-vector:nil
