module sub1 (
    in_if       if_i  , // Without modport
    int_if.mst  if_int  // With modport
);

endmodule