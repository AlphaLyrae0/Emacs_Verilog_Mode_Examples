module top (
    /*AUTOINPUT*/

    /*AUTOOUTPUT*/

);

    /*AUTOWIRE*/

    sub1 s1( /*AUTOINST*/);

    sub2 s2( /*AUTOINST*/);

endmodule
// Local Variables:
// verilog-library-flags:("-y ./sub")
// verilog-auto-inst-column:24  ;; Min. 24?
// indent-tabs-mode:nil
// End:

// verilog-auto-inst-dot-name:t
// verilog-auto-inst-vector:nil
// verilog-auto-inst-vector:nil
// verilog-auto-wire-type:"logic"
// verilog-auto-inst-sort:t
// verilog-auto-lineup:all
// verilog-auto-template-warn-unused:t
